
package CONSTANTS is
   constant IVDELAY     : time := 0 ns;
   constant NDDELAY     : time := 0 ns;
   constant NDDELAYRISE : time := 0 ns;
   constant NDDELAYFALL : time := 0 ns;
   constant NRDELAY     : time := 0 ns;
   constant DRCAS       : time := 0 ns;
   constant DRCAC       : time := 0 ns;
   constant TP_MUX      : time := 0 ns; 
   constant NumBit      : integer := 32;	
	constant NBit_Regs   : integer := 64;
	constant  NBit_addr  : integer := 5;
	   constant NBIT : integer := 32;	
end CONSTANTS;
